`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 21.02.2020 15:47:36
// Design Name: 
// Module Name: ts_muxer8
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ts_bench();
    logic [15:0] in;
    logic  [3:0]   sel;
    logic       q;
mux16 DUT(.in(in), .sel(sel), .q(q));

initial begin
//    sel = 3'b000; in = 8'b00000001; #10; //2 = 2^0 = 1
//    sel = 3'b001; in = 8'b00000010; #10; // 4 = 2^1 + 2^1
//    sel = 3'b010; in = 8'b00000100; #10; // 8 = 
//    sel = 3'b011; in = 8'b00001000; #10; // 16 = 2^4
//    sel = 3'b100; in = 8'b00010000; #10;
//    sel = 3'b101; in = 8'b00100000; #10;
//    sel = 3'b110; in = 8'b01000000; #10;
//    sel = 3'b111; in = 8'b10000000; #10;
   
//    sel = 3'b000; in = 8'b11111110; #10;
//    sel = 3'b001; in = 8'b11111101; #10;
//    sel = 3'b010; in = 8'b11111011; #10;
//    sel = 3'b011; in = 8'b11110111; #10;
//    sel = 3'b100; in = 8'b11101111; #10;
//    sel = 3'b101; in = 8'b11011111; #10;
//    sel = 3'b110; in = 8'b10111111; #10;
//    sel = 3'b111; in = 8'b01111111; #10;//2


    sel = 4'b0000; in = 16'b0000000000000001; #10; //2 = 2^0 = 1
    sel = 4'b0001; in = 16'b0000000000000010; #10; // 4 = 2^1 + 2^1
    sel = 4'b0010; in = 16'b0000000000000100; #10; // 8 = 
    sel = 4'b0011; in = 16'b0000000000001000; #10; // 16 = 2^4
    sel = 4'b0100; in = 16'b0000000000010000; #10;
    sel = 4'b0101; in = 16'b0000000000100000; #10;
    sel = 4'b0110; in = 16'b0000000001000000; #10;
    sel = 4'b0111; in = 16'b0000000010000000; #10; 
    
    sel = 4'b1000; in = 16'b0000000100000000; #10; // 4 = 2^1 + 2^1
    sel = 4'b1001; in = 16'b0000001000000000; #10; // 8 = 
    sel = 4'b1010; in = 16'b0000010000000000; #10; // 16 = 2^4
    sel = 4'b1011; in = 16'b0000100000000000; #10;
    sel = 4'b1100; in = 16'b0001000000000000; #10;
    sel = 4'b1101; in = 16'b0010000000000000; #10;
    sel = 4'b1110; in = 16'b0100000000000000; #10;
    sel = 4'b1111; in = 16'b1000000000000000; #10; //2 = 2^0 = 1

   
//    sel = 3'b000; in = 8'b11111110; #10;
//    sel = 3'b001; in = 8'b11111101; #10;
//    sel = 3'b010; in = 8'b11111011; #10;
//    sel = 3'b011; in = 8'b11110111; #10;
//    sel = 3'b100; in = 8'b11101111; #10;
//    sel = 3'b101; in = 8'b11011111; #10;
//    sel = 3'b110; in = 8'b10111111; #10;
//    sel = 3'b111; in = 8'b01111111; #10;//2^0+2
    
    
//    sel = 2'b00; in = 4'b0001; #10;
//    sel = 2'b01; in = 4'b0010; #10;
//    sel = 2'b10; in = 4'b0100; #10;
//    sel = 2'b11; in = 4'b1000; #10;
   
//    sel = 2'b00; in = 4'b1110; #10;
//    sel = 2'b01; in = 4'b1101; #10;
//    sel = 2'b10; in = 4'b1011; #10;
//    sel = 2'b11; in = 4'b0111; #10;
//  in = 0; #10
//  sel = 0; #10
//    repeat (31) begin
//        in  = (2^sel); #10;
//        sel = sel+1; #10;
//    end
//  in = 0; #10
//  sel = 0; #10
//    repeat (31) begin
//        in  = 2^32-(2^sel); #10;
//        sel = sel+1; #10;
//    end


$finish;
end;
endmodule
